package ArmFilePaths is

	--	Pfad zum Testvektorverzeichnis, betriebssystem- und und Projektabhängig;
	constant TESTVECTOR_FOLDER_PATH : STRING := "C:/HardwareLab/Blatt8/";

end package ArmFilePaths;

package body ArmFilePaths is
end package body ArmFilePaths;
